
module memory(values);
  output wire [15:0][31:0] values;



  assign values[0] = 32'b00000001100101011100000000100000;
  assign values[1] = 32'b00000000101111001010100111000000;
  assign values[2] = 32'b00000000010111001101000101100000;
  assign values[3] = 32'b00000000001011100011101000000000;
  assign values[4] = 32'b00000000000101110001011101000000;
  assign values[5] = 32'b00000000000010111000101011100000;
  assign values[6] = 32'b00000000000001011100010101100000;
  assign values[7] = 32'b00000000000000101110001010100000;
  assign values[8] = 32'b00000000000000010111000101100000;
  assign values[9] = 32'b00000000000000001011100010100000;
  assign values[10]= 32'b00000000000000000101110001100000;
  assign values[11]= 32'b00000000000000000010111000100000;
  assign values[12]= 32'b00000000000000000001011100100000;
  assign values[13]= 32'b00000000000000000000101110000000;
  assign values[14]= 32'b00000000000000000000010111000000;
  assign values[15]= 32'b00000000000000000000001011100000;

endmodule